module default_env_env;
   my_interface my_interface_inst();

   // Creating the environment components
   
   driver u_module1();
   
   monitor u_module2();
   

endmodule : default_env